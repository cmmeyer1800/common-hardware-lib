{# template/rtl/template_mod.sv #}
module {{mod_name}} #(
    // @TODO: Add Parameters Here
) (
    // @TODO: Add Ports Here
);

// @TODO: Add Logic Here
    
endmodule