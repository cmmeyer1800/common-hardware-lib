package alu_com;

typedef enum logic [2:0] { aluopADD, aluopSUB, aluopAND, aluopOR, aluopXOR, aluopSHL, aluopSHR } aluop;

endpackage